module (
    
);
    
endmodule