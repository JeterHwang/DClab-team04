module AudRecorder (
    input 


);