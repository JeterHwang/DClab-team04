module Top(
    
);
    
endmodule