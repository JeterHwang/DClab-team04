module AudPlayer (



);