module I2cIntializer(
    input i_rst_n,
    input i_clk,
    input i_start,
    output o_finished,
    output o_sclk,
    output o_sdat,
    output O_oen
);



always_comb begin
    
end

always_ff @(posedge ck, posedge arst) begin
    
end

endmodule
