module Offense_blocked_four(
    input   [4:0] X,
    input   [4:0] Y,
    input   [1:0] turn,
    output  check 
);

logic checked;

assign check = checked;

always_comb begin
    
end
endmodule