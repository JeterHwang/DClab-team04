
module SearchOffense(
    input         i_clk,
	input         i_rst_n,
	input         i_start,
	input         board i_board,         // 15*15*2 bit chess board
    input         i_turn,          
	input         i_X,
    input         i_Y,
    output        hit  
);
    
endmodule